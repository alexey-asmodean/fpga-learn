module repeater(
    input wire clk,
    output wire clk1
);

assign clk1 = clk;

endmodule